module main;
	reg [31:0] a[5:0][5:0], b[5:0][5:0]; 
	wire [31:0] result;
	calc calc0 (result,
		a[0][0],a[0][1],a[0][2],a[0][3],a[0][4],a[0][5],
		a[1][0],a[1][1],a[1][2],a[1][3],a[1][4],a[1][5],
		a[2][0],a[2][1],a[2][2],a[2][3],a[2][4],a[2][5],
		a[3][0],a[3][1],a[3][2],a[3][3],a[3][4],a[3][5],
		a[4][0],a[4][1],a[4][2],a[4][3],a[4][4],a[4][5],
		a[5][0],a[5][1],a[5][2],a[5][3],a[5][4],a[5][5],
		b[0][0],b[0][1],b[0][2],b[0][3],b[0][4],b[0][5],
		b[1][0],b[1][1],b[1][2],b[1][3],b[1][4],b[1][5],
		b[2][0],b[2][1],b[2][2],b[2][3],b[2][4],b[2][5],
		b[3][0],b[3][1],b[3][2],b[3][3],b[3][4],b[3][5],
		b[4][0],b[4][1],b[4][2],b[4][3],b[4][4],b[4][5],
		b[5][0],b[5][1],b[5][2],b[5][3],b[5][4],b[5][5]);
	
	initial
	begin
		$dumpfile("main.vcd");
		$dumpvars(0,main);
	end

	initial
	begin
		a[0][0]=3;a[0][1]=3;a[0][2]=3;a[0][3]=3;a[0][4]=3;a[0][5]=3;
		a[1][0]=3;a[1][1]=3;a[1][2]=3;a[1][3]=3;a[1][4]=3;a[1][5]=3;
		a[2][0]=3;a[2][1]=3;a[2][2]=3;a[2][3]=3;a[2][4]=3;a[2][5]=3;
		a[3][0]=3;a[3][1]=3;a[3][2]=3;a[3][3]=3;a[3][4]=3;a[3][5]=3;
		a[4][0]=3;a[4][1]=3;a[4][2]=3;a[4][3]=3;a[4][4]=3;a[4][5]=3;
		a[5][0]=3;a[5][1]=3;a[5][2]=3;a[5][3]=3;a[5][4]=3;a[5][5]=3;
		b[0][0]=3;b[0][1]=3;b[0][2]=3;b[0][3]=3;b[0][4]=3;b[0][5]=3;
		b[1][0]=3;b[1][1]=3;b[1][2]=3;b[1][3]=3;b[1][4]=3;b[1][5]=3;
		b[2][0]=3;b[2][1]=3;b[2][2]=3;b[2][3]=3;b[2][4]=3;b[2][5]=3;
		b[3][0]=3;b[3][1]=3;b[3][2]=3;b[3][3]=3;b[3][4]=3;b[3][5]=3;
		b[4][0]=3;b[4][1]=3;b[4][2]=3;b[4][3]=3;b[4][4]=3;b[4][5]=3;
		b[5][0]=3;b[5][1]=3;b[5][2]=3;b[5][3]=3;b[5][4]=3;b[5][5]=3;
		#1 $stop;
		end

endmodule
