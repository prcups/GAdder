module main;
	reg [31:0] a[5:0][5:0], b[5:0][5:0];
	reg [31:0] result;
	reg [7:0] i, j;

	initial
		begin
			$dumpfile("main.vcd");
			$dumpvars(0,main);
		end
		
		initial
		begin
			a[0][0]=3;a[0][1]=3;a[0][2]=3;a[0][3]=3;a[0][4]=3;a[0][5]=3;
			a[1][0]=3;a[1][1]=3;a[1][2]=3;a[1][3]=3;a[1][4]=3;a[1][5]=3;
			a[2][0]=3;a[2][1]=3;a[2][2]=3;a[2][3]=3;a[2][4]=3;a[2][5]=3;
			a[3][0]=3;a[3][1]=3;a[3][2]=3;a[3][3]=3;a[3][4]=3;a[3][5]=3;
			a[4][0]=3;a[4][1]=3;a[4][2]=3;a[4][3]=3;a[4][4]=3;a[4][5]=3;
			a[5][0]=3;a[5][1]=3;a[5][2]=3;a[5][3]=3;a[5][4]=3;a[5][5]=3;
			
			b[0][0]=3;b[0][1]=3;b[0][2]=3;b[0][3]=3;b[0][4]=3;b[0][5]=3;
			b[1][0]=3;b[1][1]=3;b[1][2]=3;b[1][3]=3;b[1][4]=3;b[1][5]=3;
			b[2][0]=3;b[2][1]=3;b[2][2]=3;b[2][3]=3;b[2][4]=3;b[2][5]=3;
			b[3][0]=3;b[3][1]=3;b[3][2]=3;b[3][3]=3;b[3][4]=3;b[3][5]=3;
			b[4][0]=3;b[4][1]=3;b[4][2]=3;b[4][3]=3;b[4][4]=3;b[4][5]=3;
			b[5][0]=3;b[5][1]=3;b[5][2]=3;b[5][3]=3;b[5][4]=3;b[5][5]=3;
			
			result = 0;
			for (i = 0; i <= 5; i = i + 1)
			begin
				for (j = 0; j <= 5; j = j + 1)
				begin
				result = result + a[i][j] * b[i][j];
				end
			end
			#5 $stop;
		end

endmodule

