module multiply(F, X1, X2);
	input [31:0] X1, X2;
	output [31:0] F;
	wire [31:0] PT, T, P;
	
	buf(PT[31], 1'b0);
	buf(PT[30], 1'b0);
	buf(PT[29], 1'b0);
	buf(PT[28], 1'b0);
	buf(PT[27], 1'b0);
	buf(PT[26], 1'b0);
	buf(PT[25], 1'b0);
	buf(PT[24], 1'b0);
	buf(PT[23], 1'b0);
	buf(PT[22], 1'b0);
	buf(PT[21], 1'b0);
	buf(PT[20], 1'b0);
	buf(PT[19], 1'b0);
	buf(PT[18], 1'b0);
	buf(PT[17], 1'b0);
	buf(PT[16], 1'b0);
	buf(PT[15], 1'b0);
	buf(PT[14], 1'b0);
	buf(PT[13], 1'b0);
	buf(PT[12], 1'b0);
	buf(PT[11], 1'b0);
	buf(PT[10], 1'b0);
	buf(PT[9], 1'b0);
	buf(PT[8], 1'b0);
	buf(PT[7], 1'b0);
	buf(PT[6], 1'b0);
	buf(PT[5], 1'b0);
	buf(PT[4], 1'b0);
	buf(PT[3], 1'b0);
	buf(PT[2], 1'b0);
	buf(PT[1], 1'b0);
	buf(PT[0], 1'b0);
	and(P[31], X1[31], X2[31]);
	and(P[30], X1[30], X2[31]);
	and(P[29], X1[29], X2[31]);
	and(P[28], X1[28], X2[31]);
	and(P[27], X1[27], X2[31]);
	and(P[26], X1[26], X2[31]);
	and(P[25], X1[25], X2[31]);
	and(P[24], X1[24], X2[31]);
	and(P[23], X1[23], X2[31]);
	and(P[22], X1[22], X2[31]);
	and(P[21], X1[21], X2[31]);
	and(P[20], X1[20], X2[31]);
	and(P[19], X1[19], X2[31]);
	and(P[18], X1[18], X2[31]);
	and(P[17], X1[17], X2[31]);
	and(P[16], X1[16], X2[31]);
	and(P[15], X1[15], X2[31]);
	and(P[14], X1[14], X2[31]);
	and(P[13], X1[13], X2[31]);
	and(P[12], X1[12], X2[31]);
	and(P[11], X1[11], X2[31]);
	and(P[10], X1[10], X2[31]);
	and(P[9], X1[9], X2[31]);
	and(P[8], X1[8], X2[31]);
	and(P[7], X1[7], X2[31]);
	and(P[6], X1[6], X2[31]);
	and(P[5], X1[5], X2[31]);
	and(P[4], X1[4], X2[31]);
	and(P[3], X1[3], X2[31]);
	and(P[2], X1[2], X2[31]);
	and(P[1], X1[1], X2[31]);
	and(P[0], X1[0], X2[31]);
	fulladd fadd31 (T, PT, P);
	leftmove lm31 (PT, T);
	and(P[31], X1[31], X2[30]);
	and(P[30], X1[30], X2[30]);
	and(P[29], X1[29], X2[30]);
	and(P[28], X1[28], X2[30]);
	and(P[27], X1[27], X2[30]);
	and(P[26], X1[26], X2[30]);
	and(P[25], X1[25], X2[30]);
	and(P[24], X1[24], X2[30]);
	and(P[23], X1[23], X2[30]);
	and(P[22], X1[22], X2[30]);
	and(P[21], X1[21], X2[30]);
	and(P[20], X1[20], X2[30]);
	and(P[19], X1[19], X2[30]);
	and(P[18], X1[18], X2[30]);
	and(P[17], X1[17], X2[30]);
	and(P[16], X1[16], X2[30]);
	and(P[15], X1[15], X2[30]);
	and(P[14], X1[14], X2[30]);
	and(P[13], X1[13], X2[30]);
	and(P[12], X1[12], X2[30]);
	and(P[11], X1[11], X2[30]);
	and(P[10], X1[10], X2[30]);
	and(P[9], X1[9], X2[30]);
	and(P[8], X1[8], X2[30]);
	and(P[7], X1[7], X2[30]);
	and(P[6], X1[6], X2[30]);
	and(P[5], X1[5], X2[30]);
	and(P[4], X1[4], X2[30]);
	and(P[3], X1[3], X2[30]);
	and(P[2], X1[2], X2[30]);
	and(P[1], X1[1], X2[30]);
	and(P[0], X1[0], X2[30]);
	fulladd fadd30 (T, PT, P);
	leftmove lm30 (PT, T);
	and(P[31], X1[31], X2[29]);
	and(P[30], X1[30], X2[29]);
	and(P[29], X1[29], X2[29]);
	and(P[28], X1[28], X2[29]);
	and(P[27], X1[27], X2[29]);
	and(P[26], X1[26], X2[29]);
	and(P[25], X1[25], X2[29]);
	and(P[24], X1[24], X2[29]);
	and(P[23], X1[23], X2[29]);
	and(P[22], X1[22], X2[29]);
	and(P[21], X1[21], X2[29]);
	and(P[20], X1[20], X2[29]);
	and(P[19], X1[19], X2[29]);
	and(P[18], X1[18], X2[29]);
	and(P[17], X1[17], X2[29]);
	and(P[16], X1[16], X2[29]);
	and(P[15], X1[15], X2[29]);
	and(P[14], X1[14], X2[29]);
	and(P[13], X1[13], X2[29]);
	and(P[12], X1[12], X2[29]);
	and(P[11], X1[11], X2[29]);
	and(P[10], X1[10], X2[29]);
	and(P[9], X1[9], X2[29]);
	and(P[8], X1[8], X2[29]);
	and(P[7], X1[7], X2[29]);
	and(P[6], X1[6], X2[29]);
	and(P[5], X1[5], X2[29]);
	and(P[4], X1[4], X2[29]);
	and(P[3], X1[3], X2[29]);
	and(P[2], X1[2], X2[29]);
	and(P[1], X1[1], X2[29]);
	and(P[0], X1[0], X2[29]);
	fulladd fadd29 (T, PT, P);
	leftmove lm29 (PT, T);
	and(P[31], X1[31], X2[28]);
	and(P[30], X1[30], X2[28]);
	and(P[29], X1[29], X2[28]);
	and(P[28], X1[28], X2[28]);
	and(P[27], X1[27], X2[28]);
	and(P[26], X1[26], X2[28]);
	and(P[25], X1[25], X2[28]);
	and(P[24], X1[24], X2[28]);
	and(P[23], X1[23], X2[28]);
	and(P[22], X1[22], X2[28]);
	and(P[21], X1[21], X2[28]);
	and(P[20], X1[20], X2[28]);
	and(P[19], X1[19], X2[28]);
	and(P[18], X1[18], X2[28]);
	and(P[17], X1[17], X2[28]);
	and(P[16], X1[16], X2[28]);
	and(P[15], X1[15], X2[28]);
	and(P[14], X1[14], X2[28]);
	and(P[13], X1[13], X2[28]);
	and(P[12], X1[12], X2[28]);
	and(P[11], X1[11], X2[28]);
	and(P[10], X1[10], X2[28]);
	and(P[9], X1[9], X2[28]);
	and(P[8], X1[8], X2[28]);
	and(P[7], X1[7], X2[28]);
	and(P[6], X1[6], X2[28]);
	and(P[5], X1[5], X2[28]);
	and(P[4], X1[4], X2[28]);
	and(P[3], X1[3], X2[28]);
	and(P[2], X1[2], X2[28]);
	and(P[1], X1[1], X2[28]);
	and(P[0], X1[0], X2[28]);
	fulladd fadd28 (T, PT, P);
	leftmove lm28 (PT, T);
	and(P[31], X1[31], X2[27]);
	and(P[30], X1[30], X2[27]);
	and(P[29], X1[29], X2[27]);
	and(P[28], X1[28], X2[27]);
	and(P[27], X1[27], X2[27]);
	and(P[26], X1[26], X2[27]);
	and(P[25], X1[25], X2[27]);
	and(P[24], X1[24], X2[27]);
	and(P[23], X1[23], X2[27]);
	and(P[22], X1[22], X2[27]);
	and(P[21], X1[21], X2[27]);
	and(P[20], X1[20], X2[27]);
	and(P[19], X1[19], X2[27]);
	and(P[18], X1[18], X2[27]);
	and(P[17], X1[17], X2[27]);
	and(P[16], X1[16], X2[27]);
	and(P[15], X1[15], X2[27]);
	and(P[14], X1[14], X2[27]);
	and(P[13], X1[13], X2[27]);
	and(P[12], X1[12], X2[27]);
	and(P[11], X1[11], X2[27]);
	and(P[10], X1[10], X2[27]);
	and(P[9], X1[9], X2[27]);
	and(P[8], X1[8], X2[27]);
	and(P[7], X1[7], X2[27]);
	and(P[6], X1[6], X2[27]);
	and(P[5], X1[5], X2[27]);
	and(P[4], X1[4], X2[27]);
	and(P[3], X1[3], X2[27]);
	and(P[2], X1[2], X2[27]);
	and(P[1], X1[1], X2[27]);
	and(P[0], X1[0], X2[27]);
	fulladd fadd27 (T, PT, P);
	leftmove lm27 (PT, T);
	and(P[31], X1[31], X2[26]);
	and(P[30], X1[30], X2[26]);
	and(P[29], X1[29], X2[26]);
	and(P[28], X1[28], X2[26]);
	and(P[27], X1[27], X2[26]);
	and(P[26], X1[26], X2[26]);
	and(P[25], X1[25], X2[26]);
	and(P[24], X1[24], X2[26]);
	and(P[23], X1[23], X2[26]);
	and(P[22], X1[22], X2[26]);
	and(P[21], X1[21], X2[26]);
	and(P[20], X1[20], X2[26]);
	and(P[19], X1[19], X2[26]);
	and(P[18], X1[18], X2[26]);
	and(P[17], X1[17], X2[26]);
	and(P[16], X1[16], X2[26]);
	and(P[15], X1[15], X2[26]);
	and(P[14], X1[14], X2[26]);
	and(P[13], X1[13], X2[26]);
	and(P[12], X1[12], X2[26]);
	and(P[11], X1[11], X2[26]);
	and(P[10], X1[10], X2[26]);
	and(P[9], X1[9], X2[26]);
	and(P[8], X1[8], X2[26]);
	and(P[7], X1[7], X2[26]);
	and(P[6], X1[6], X2[26]);
	and(P[5], X1[5], X2[26]);
	and(P[4], X1[4], X2[26]);
	and(P[3], X1[3], X2[26]);
	and(P[2], X1[2], X2[26]);
	and(P[1], X1[1], X2[26]);
	and(P[0], X1[0], X2[26]);
	fulladd fadd26 (T, PT, P);
	leftmove lm26 (PT, T);
	and(P[31], X1[31], X2[25]);
	and(P[30], X1[30], X2[25]);
	and(P[29], X1[29], X2[25]);
	and(P[28], X1[28], X2[25]);
	and(P[27], X1[27], X2[25]);
	and(P[26], X1[26], X2[25]);
	and(P[25], X1[25], X2[25]);
	and(P[24], X1[24], X2[25]);
	and(P[23], X1[23], X2[25]);
	and(P[22], X1[22], X2[25]);
	and(P[21], X1[21], X2[25]);
	and(P[20], X1[20], X2[25]);
	and(P[19], X1[19], X2[25]);
	and(P[18], X1[18], X2[25]);
	and(P[17], X1[17], X2[25]);
	and(P[16], X1[16], X2[25]);
	and(P[15], X1[15], X2[25]);
	and(P[14], X1[14], X2[25]);
	and(P[13], X1[13], X2[25]);
	and(P[12], X1[12], X2[25]);
	and(P[11], X1[11], X2[25]);
	and(P[10], X1[10], X2[25]);
	and(P[9], X1[9], X2[25]);
	and(P[8], X1[8], X2[25]);
	and(P[7], X1[7], X2[25]);
	and(P[6], X1[6], X2[25]);
	and(P[5], X1[5], X2[25]);
	and(P[4], X1[4], X2[25]);
	and(P[3], X1[3], X2[25]);
	and(P[2], X1[2], X2[25]);
	and(P[1], X1[1], X2[25]);
	and(P[0], X1[0], X2[25]);
	fulladd fadd25 (T, PT, P);
	leftmove lm25 (PT, T);
	and(P[31], X1[31], X2[24]);
	and(P[30], X1[30], X2[24]);
	and(P[29], X1[29], X2[24]);
	and(P[28], X1[28], X2[24]);
	and(P[27], X1[27], X2[24]);
	and(P[26], X1[26], X2[24]);
	and(P[25], X1[25], X2[24]);
	and(P[24], X1[24], X2[24]);
	and(P[23], X1[23], X2[24]);
	and(P[22], X1[22], X2[24]);
	and(P[21], X1[21], X2[24]);
	and(P[20], X1[20], X2[24]);
	and(P[19], X1[19], X2[24]);
	and(P[18], X1[18], X2[24]);
	and(P[17], X1[17], X2[24]);
	and(P[16], X1[16], X2[24]);
	and(P[15], X1[15], X2[24]);
	and(P[14], X1[14], X2[24]);
	and(P[13], X1[13], X2[24]);
	and(P[12], X1[12], X2[24]);
	and(P[11], X1[11], X2[24]);
	and(P[10], X1[10], X2[24]);
	and(P[9], X1[9], X2[24]);
	and(P[8], X1[8], X2[24]);
	and(P[7], X1[7], X2[24]);
	and(P[6], X1[6], X2[24]);
	and(P[5], X1[5], X2[24]);
	and(P[4], X1[4], X2[24]);
	and(P[3], X1[3], X2[24]);
	and(P[2], X1[2], X2[24]);
	and(P[1], X1[1], X2[24]);
	and(P[0], X1[0], X2[24]);
	fulladd fadd24 (T, PT, P);
	leftmove lm24 (PT, T);
	and(P[31], X1[31], X2[23]);
	and(P[30], X1[30], X2[23]);
	and(P[29], X1[29], X2[23]);
	and(P[28], X1[28], X2[23]);
	and(P[27], X1[27], X2[23]);
	and(P[26], X1[26], X2[23]);
	and(P[25], X1[25], X2[23]);
	and(P[24], X1[24], X2[23]);
	and(P[23], X1[23], X2[23]);
	and(P[22], X1[22], X2[23]);
	and(P[21], X1[21], X2[23]);
	and(P[20], X1[20], X2[23]);
	and(P[19], X1[19], X2[23]);
	and(P[18], X1[18], X2[23]);
	and(P[17], X1[17], X2[23]);
	and(P[16], X1[16], X2[23]);
	and(P[15], X1[15], X2[23]);
	and(P[14], X1[14], X2[23]);
	and(P[13], X1[13], X2[23]);
	and(P[12], X1[12], X2[23]);
	and(P[11], X1[11], X2[23]);
	and(P[10], X1[10], X2[23]);
	and(P[9], X1[9], X2[23]);
	and(P[8], X1[8], X2[23]);
	and(P[7], X1[7], X2[23]);
	and(P[6], X1[6], X2[23]);
	and(P[5], X1[5], X2[23]);
	and(P[4], X1[4], X2[23]);
	and(P[3], X1[3], X2[23]);
	and(P[2], X1[2], X2[23]);
	and(P[1], X1[1], X2[23]);
	and(P[0], X1[0], X2[23]);
	fulladd fadd23 (T, PT, P);
	leftmove lm23 (PT, T);
	and(P[31], X1[31], X2[22]);
	and(P[30], X1[30], X2[22]);
	and(P[29], X1[29], X2[22]);
	and(P[28], X1[28], X2[22]);
	and(P[27], X1[27], X2[22]);
	and(P[26], X1[26], X2[22]);
	and(P[25], X1[25], X2[22]);
	and(P[24], X1[24], X2[22]);
	and(P[23], X1[23], X2[22]);
	and(P[22], X1[22], X2[22]);
	and(P[21], X1[21], X2[22]);
	and(P[20], X1[20], X2[22]);
	and(P[19], X1[19], X2[22]);
	and(P[18], X1[18], X2[22]);
	and(P[17], X1[17], X2[22]);
	and(P[16], X1[16], X2[22]);
	and(P[15], X1[15], X2[22]);
	and(P[14], X1[14], X2[22]);
	and(P[13], X1[13], X2[22]);
	and(P[12], X1[12], X2[22]);
	and(P[11], X1[11], X2[22]);
	and(P[10], X1[10], X2[22]);
	and(P[9], X1[9], X2[22]);
	and(P[8], X1[8], X2[22]);
	and(P[7], X1[7], X2[22]);
	and(P[6], X1[6], X2[22]);
	and(P[5], X1[5], X2[22]);
	and(P[4], X1[4], X2[22]);
	and(P[3], X1[3], X2[22]);
	and(P[2], X1[2], X2[22]);
	and(P[1], X1[1], X2[22]);
	and(P[0], X1[0], X2[22]);
	fulladd fadd22 (T, PT, P);
	leftmove lm22 (PT, T);
	and(P[31], X1[31], X2[21]);
	and(P[30], X1[30], X2[21]);
	and(P[29], X1[29], X2[21]);
	and(P[28], X1[28], X2[21]);
	and(P[27], X1[27], X2[21]);
	and(P[26], X1[26], X2[21]);
	and(P[25], X1[25], X2[21]);
	and(P[24], X1[24], X2[21]);
	and(P[23], X1[23], X2[21]);
	and(P[22], X1[22], X2[21]);
	and(P[21], X1[21], X2[21]);
	and(P[20], X1[20], X2[21]);
	and(P[19], X1[19], X2[21]);
	and(P[18], X1[18], X2[21]);
	and(P[17], X1[17], X2[21]);
	and(P[16], X1[16], X2[21]);
	and(P[15], X1[15], X2[21]);
	and(P[14], X1[14], X2[21]);
	and(P[13], X1[13], X2[21]);
	and(P[12], X1[12], X2[21]);
	and(P[11], X1[11], X2[21]);
	and(P[10], X1[10], X2[21]);
	and(P[9], X1[9], X2[21]);
	and(P[8], X1[8], X2[21]);
	and(P[7], X1[7], X2[21]);
	and(P[6], X1[6], X2[21]);
	and(P[5], X1[5], X2[21]);
	and(P[4], X1[4], X2[21]);
	and(P[3], X1[3], X2[21]);
	and(P[2], X1[2], X2[21]);
	and(P[1], X1[1], X2[21]);
	and(P[0], X1[0], X2[21]);
	fulladd fadd21 (T, PT, P);
	leftmove lm21 (PT, T);
	and(P[31], X1[31], X2[20]);
	and(P[30], X1[30], X2[20]);
	and(P[29], X1[29], X2[20]);
	and(P[28], X1[28], X2[20]);
	and(P[27], X1[27], X2[20]);
	and(P[26], X1[26], X2[20]);
	and(P[25], X1[25], X2[20]);
	and(P[24], X1[24], X2[20]);
	and(P[23], X1[23], X2[20]);
	and(P[22], X1[22], X2[20]);
	and(P[21], X1[21], X2[20]);
	and(P[20], X1[20], X2[20]);
	and(P[19], X1[19], X2[20]);
	and(P[18], X1[18], X2[20]);
	and(P[17], X1[17], X2[20]);
	and(P[16], X1[16], X2[20]);
	and(P[15], X1[15], X2[20]);
	and(P[14], X1[14], X2[20]);
	and(P[13], X1[13], X2[20]);
	and(P[12], X1[12], X2[20]);
	and(P[11], X1[11], X2[20]);
	and(P[10], X1[10], X2[20]);
	and(P[9], X1[9], X2[20]);
	and(P[8], X1[8], X2[20]);
	and(P[7], X1[7], X2[20]);
	and(P[6], X1[6], X2[20]);
	and(P[5], X1[5], X2[20]);
	and(P[4], X1[4], X2[20]);
	and(P[3], X1[3], X2[20]);
	and(P[2], X1[2], X2[20]);
	and(P[1], X1[1], X2[20]);
	and(P[0], X1[0], X2[20]);
	fulladd fadd20 (T, PT, P);
	leftmove lm20 (PT, T);
	and(P[31], X1[31], X2[19]);
	and(P[30], X1[30], X2[19]);
	and(P[29], X1[29], X2[19]);
	and(P[28], X1[28], X2[19]);
	and(P[27], X1[27], X2[19]);
	and(P[26], X1[26], X2[19]);
	and(P[25], X1[25], X2[19]);
	and(P[24], X1[24], X2[19]);
	and(P[23], X1[23], X2[19]);
	and(P[22], X1[22], X2[19]);
	and(P[21], X1[21], X2[19]);
	and(P[20], X1[20], X2[19]);
	and(P[19], X1[19], X2[19]);
	and(P[18], X1[18], X2[19]);
	and(P[17], X1[17], X2[19]);
	and(P[16], X1[16], X2[19]);
	and(P[15], X1[15], X2[19]);
	and(P[14], X1[14], X2[19]);
	and(P[13], X1[13], X2[19]);
	and(P[12], X1[12], X2[19]);
	and(P[11], X1[11], X2[19]);
	and(P[10], X1[10], X2[19]);
	and(P[9], X1[9], X2[19]);
	and(P[8], X1[8], X2[19]);
	and(P[7], X1[7], X2[19]);
	and(P[6], X1[6], X2[19]);
	and(P[5], X1[5], X2[19]);
	and(P[4], X1[4], X2[19]);
	and(P[3], X1[3], X2[19]);
	and(P[2], X1[2], X2[19]);
	and(P[1], X1[1], X2[19]);
	and(P[0], X1[0], X2[19]);
	fulladd fadd19 (T, PT, P);
	leftmove lm19 (PT, T);
	and(P[31], X1[31], X2[18]);
	and(P[30], X1[30], X2[18]);
	and(P[29], X1[29], X2[18]);
	and(P[28], X1[28], X2[18]);
	and(P[27], X1[27], X2[18]);
	and(P[26], X1[26], X2[18]);
	and(P[25], X1[25], X2[18]);
	and(P[24], X1[24], X2[18]);
	and(P[23], X1[23], X2[18]);
	and(P[22], X1[22], X2[18]);
	and(P[21], X1[21], X2[18]);
	and(P[20], X1[20], X2[18]);
	and(P[19], X1[19], X2[18]);
	and(P[18], X1[18], X2[18]);
	and(P[17], X1[17], X2[18]);
	and(P[16], X1[16], X2[18]);
	and(P[15], X1[15], X2[18]);
	and(P[14], X1[14], X2[18]);
	and(P[13], X1[13], X2[18]);
	and(P[12], X1[12], X2[18]);
	and(P[11], X1[11], X2[18]);
	and(P[10], X1[10], X2[18]);
	and(P[9], X1[9], X2[18]);
	and(P[8], X1[8], X2[18]);
	and(P[7], X1[7], X2[18]);
	and(P[6], X1[6], X2[18]);
	and(P[5], X1[5], X2[18]);
	and(P[4], X1[4], X2[18]);
	and(P[3], X1[3], X2[18]);
	and(P[2], X1[2], X2[18]);
	and(P[1], X1[1], X2[18]);
	and(P[0], X1[0], X2[18]);
	fulladd fadd18 (T, PT, P);
	leftmove lm18 (PT, T);
	and(P[31], X1[31], X2[17]);
	and(P[30], X1[30], X2[17]);
	and(P[29], X1[29], X2[17]);
	and(P[28], X1[28], X2[17]);
	and(P[27], X1[27], X2[17]);
	and(P[26], X1[26], X2[17]);
	and(P[25], X1[25], X2[17]);
	and(P[24], X1[24], X2[17]);
	and(P[23], X1[23], X2[17]);
	and(P[22], X1[22], X2[17]);
	and(P[21], X1[21], X2[17]);
	and(P[20], X1[20], X2[17]);
	and(P[19], X1[19], X2[17]);
	and(P[18], X1[18], X2[17]);
	and(P[17], X1[17], X2[17]);
	and(P[16], X1[16], X2[17]);
	and(P[15], X1[15], X2[17]);
	and(P[14], X1[14], X2[17]);
	and(P[13], X1[13], X2[17]);
	and(P[12], X1[12], X2[17]);
	and(P[11], X1[11], X2[17]);
	and(P[10], X1[10], X2[17]);
	and(P[9], X1[9], X2[17]);
	and(P[8], X1[8], X2[17]);
	and(P[7], X1[7], X2[17]);
	and(P[6], X1[6], X2[17]);
	and(P[5], X1[5], X2[17]);
	and(P[4], X1[4], X2[17]);
	and(P[3], X1[3], X2[17]);
	and(P[2], X1[2], X2[17]);
	and(P[1], X1[1], X2[17]);
	and(P[0], X1[0], X2[17]);
	fulladd fadd17 (T, PT, P);
	leftmove lm17 (PT, T);
	and(P[31], X1[31], X2[16]);
	and(P[30], X1[30], X2[16]);
	and(P[29], X1[29], X2[16]);
	and(P[28], X1[28], X2[16]);
	and(P[27], X1[27], X2[16]);
	and(P[26], X1[26], X2[16]);
	and(P[25], X1[25], X2[16]);
	and(P[24], X1[24], X2[16]);
	and(P[23], X1[23], X2[16]);
	and(P[22], X1[22], X2[16]);
	and(P[21], X1[21], X2[16]);
	and(P[20], X1[20], X2[16]);
	and(P[19], X1[19], X2[16]);
	and(P[18], X1[18], X2[16]);
	and(P[17], X1[17], X2[16]);
	and(P[16], X1[16], X2[16]);
	and(P[15], X1[15], X2[16]);
	and(P[14], X1[14], X2[16]);
	and(P[13], X1[13], X2[16]);
	and(P[12], X1[12], X2[16]);
	and(P[11], X1[11], X2[16]);
	and(P[10], X1[10], X2[16]);
	and(P[9], X1[9], X2[16]);
	and(P[8], X1[8], X2[16]);
	and(P[7], X1[7], X2[16]);
	and(P[6], X1[6], X2[16]);
	and(P[5], X1[5], X2[16]);
	and(P[4], X1[4], X2[16]);
	and(P[3], X1[3], X2[16]);
	and(P[2], X1[2], X2[16]);
	and(P[1], X1[1], X2[16]);
	and(P[0], X1[0], X2[16]);
	fulladd fadd16 (T, PT, P);
	leftmove lm16 (PT, T);
	and(P[31], X1[31], X2[15]);
	and(P[30], X1[30], X2[15]);
	and(P[29], X1[29], X2[15]);
	and(P[28], X1[28], X2[15]);
	and(P[27], X1[27], X2[15]);
	and(P[26], X1[26], X2[15]);
	and(P[25], X1[25], X2[15]);
	and(P[24], X1[24], X2[15]);
	and(P[23], X1[23], X2[15]);
	and(P[22], X1[22], X2[15]);
	and(P[21], X1[21], X2[15]);
	and(P[20], X1[20], X2[15]);
	and(P[19], X1[19], X2[15]);
	and(P[18], X1[18], X2[15]);
	and(P[17], X1[17], X2[15]);
	and(P[16], X1[16], X2[15]);
	and(P[15], X1[15], X2[15]);
	and(P[14], X1[14], X2[15]);
	and(P[13], X1[13], X2[15]);
	and(P[12], X1[12], X2[15]);
	and(P[11], X1[11], X2[15]);
	and(P[10], X1[10], X2[15]);
	and(P[9], X1[9], X2[15]);
	and(P[8], X1[8], X2[15]);
	and(P[7], X1[7], X2[15]);
	and(P[6], X1[6], X2[15]);
	and(P[5], X1[5], X2[15]);
	and(P[4], X1[4], X2[15]);
	and(P[3], X1[3], X2[15]);
	and(P[2], X1[2], X2[15]);
	and(P[1], X1[1], X2[15]);
	and(P[0], X1[0], X2[15]);
	fulladd fadd15 (T, PT, P);
	leftmove lm15 (PT, T);
	and(P[31], X1[31], X2[14]);
	and(P[30], X1[30], X2[14]);
	and(P[29], X1[29], X2[14]);
	and(P[28], X1[28], X2[14]);
	and(P[27], X1[27], X2[14]);
	and(P[26], X1[26], X2[14]);
	and(P[25], X1[25], X2[14]);
	and(P[24], X1[24], X2[14]);
	and(P[23], X1[23], X2[14]);
	and(P[22], X1[22], X2[14]);
	and(P[21], X1[21], X2[14]);
	and(P[20], X1[20], X2[14]);
	and(P[19], X1[19], X2[14]);
	and(P[18], X1[18], X2[14]);
	and(P[17], X1[17], X2[14]);
	and(P[16], X1[16], X2[14]);
	and(P[15], X1[15], X2[14]);
	and(P[14], X1[14], X2[14]);
	and(P[13], X1[13], X2[14]);
	and(P[12], X1[12], X2[14]);
	and(P[11], X1[11], X2[14]);
	and(P[10], X1[10], X2[14]);
	and(P[9], X1[9], X2[14]);
	and(P[8], X1[8], X2[14]);
	and(P[7], X1[7], X2[14]);
	and(P[6], X1[6], X2[14]);
	and(P[5], X1[5], X2[14]);
	and(P[4], X1[4], X2[14]);
	and(P[3], X1[3], X2[14]);
	and(P[2], X1[2], X2[14]);
	and(P[1], X1[1], X2[14]);
	and(P[0], X1[0], X2[14]);
	fulladd fadd14 (T, PT, P);
	leftmove lm14 (PT, T);
	and(P[31], X1[31], X2[13]);
	and(P[30], X1[30], X2[13]);
	and(P[29], X1[29], X2[13]);
	and(P[28], X1[28], X2[13]);
	and(P[27], X1[27], X2[13]);
	and(P[26], X1[26], X2[13]);
	and(P[25], X1[25], X2[13]);
	and(P[24], X1[24], X2[13]);
	and(P[23], X1[23], X2[13]);
	and(P[22], X1[22], X2[13]);
	and(P[21], X1[21], X2[13]);
	and(P[20], X1[20], X2[13]);
	and(P[19], X1[19], X2[13]);
	and(P[18], X1[18], X2[13]);
	and(P[17], X1[17], X2[13]);
	and(P[16], X1[16], X2[13]);
	and(P[15], X1[15], X2[13]);
	and(P[14], X1[14], X2[13]);
	and(P[13], X1[13], X2[13]);
	and(P[12], X1[12], X2[13]);
	and(P[11], X1[11], X2[13]);
	and(P[10], X1[10], X2[13]);
	and(P[9], X1[9], X2[13]);
	and(P[8], X1[8], X2[13]);
	and(P[7], X1[7], X2[13]);
	and(P[6], X1[6], X2[13]);
	and(P[5], X1[5], X2[13]);
	and(P[4], X1[4], X2[13]);
	and(P[3], X1[3], X2[13]);
	and(P[2], X1[2], X2[13]);
	and(P[1], X1[1], X2[13]);
	and(P[0], X1[0], X2[13]);
	fulladd fadd13 (T, PT, P);
	leftmove lm13 (PT, T);
	and(P[31], X1[31], X2[12]);
	and(P[30], X1[30], X2[12]);
	and(P[29], X1[29], X2[12]);
	and(P[28], X1[28], X2[12]);
	and(P[27], X1[27], X2[12]);
	and(P[26], X1[26], X2[12]);
	and(P[25], X1[25], X2[12]);
	and(P[24], X1[24], X2[12]);
	and(P[23], X1[23], X2[12]);
	and(P[22], X1[22], X2[12]);
	and(P[21], X1[21], X2[12]);
	and(P[20], X1[20], X2[12]);
	and(P[19], X1[19], X2[12]);
	and(P[18], X1[18], X2[12]);
	and(P[17], X1[17], X2[12]);
	and(P[16], X1[16], X2[12]);
	and(P[15], X1[15], X2[12]);
	and(P[14], X1[14], X2[12]);
	and(P[13], X1[13], X2[12]);
	and(P[12], X1[12], X2[12]);
	and(P[11], X1[11], X2[12]);
	and(P[10], X1[10], X2[12]);
	and(P[9], X1[9], X2[12]);
	and(P[8], X1[8], X2[12]);
	and(P[7], X1[7], X2[12]);
	and(P[6], X1[6], X2[12]);
	and(P[5], X1[5], X2[12]);
	and(P[4], X1[4], X2[12]);
	and(P[3], X1[3], X2[12]);
	and(P[2], X1[2], X2[12]);
	and(P[1], X1[1], X2[12]);
	and(P[0], X1[0], X2[12]);
	fulladd fadd12 (T, PT, P);
	leftmove lm12 (PT, T);
	and(P[31], X1[31], X2[11]);
	and(P[30], X1[30], X2[11]);
	and(P[29], X1[29], X2[11]);
	and(P[28], X1[28], X2[11]);
	and(P[27], X1[27], X2[11]);
	and(P[26], X1[26], X2[11]);
	and(P[25], X1[25], X2[11]);
	and(P[24], X1[24], X2[11]);
	and(P[23], X1[23], X2[11]);
	and(P[22], X1[22], X2[11]);
	and(P[21], X1[21], X2[11]);
	and(P[20], X1[20], X2[11]);
	and(P[19], X1[19], X2[11]);
	and(P[18], X1[18], X2[11]);
	and(P[17], X1[17], X2[11]);
	and(P[16], X1[16], X2[11]);
	and(P[15], X1[15], X2[11]);
	and(P[14], X1[14], X2[11]);
	and(P[13], X1[13], X2[11]);
	and(P[12], X1[12], X2[11]);
	and(P[11], X1[11], X2[11]);
	and(P[10], X1[10], X2[11]);
	and(P[9], X1[9], X2[11]);
	and(P[8], X1[8], X2[11]);
	and(P[7], X1[7], X2[11]);
	and(P[6], X1[6], X2[11]);
	and(P[5], X1[5], X2[11]);
	and(P[4], X1[4], X2[11]);
	and(P[3], X1[3], X2[11]);
	and(P[2], X1[2], X2[11]);
	and(P[1], X1[1], X2[11]);
	and(P[0], X1[0], X2[11]);
	fulladd fadd11 (T, PT, P);
	leftmove lm11 (PT, T);
	and(P[31], X1[31], X2[10]);
	and(P[30], X1[30], X2[10]);
	and(P[29], X1[29], X2[10]);
	and(P[28], X1[28], X2[10]);
	and(P[27], X1[27], X2[10]);
	and(P[26], X1[26], X2[10]);
	and(P[25], X1[25], X2[10]);
	and(P[24], X1[24], X2[10]);
	and(P[23], X1[23], X2[10]);
	and(P[22], X1[22], X2[10]);
	and(P[21], X1[21], X2[10]);
	and(P[20], X1[20], X2[10]);
	and(P[19], X1[19], X2[10]);
	and(P[18], X1[18], X2[10]);
	and(P[17], X1[17], X2[10]);
	and(P[16], X1[16], X2[10]);
	and(P[15], X1[15], X2[10]);
	and(P[14], X1[14], X2[10]);
	and(P[13], X1[13], X2[10]);
	and(P[12], X1[12], X2[10]);
	and(P[11], X1[11], X2[10]);
	and(P[10], X1[10], X2[10]);
	and(P[9], X1[9], X2[10]);
	and(P[8], X1[8], X2[10]);
	and(P[7], X1[7], X2[10]);
	and(P[6], X1[6], X2[10]);
	and(P[5], X1[5], X2[10]);
	and(P[4], X1[4], X2[10]);
	and(P[3], X1[3], X2[10]);
	and(P[2], X1[2], X2[10]);
	and(P[1], X1[1], X2[10]);
	and(P[0], X1[0], X2[10]);
	fulladd fadd10 (T, PT, P);
	leftmove lm10 (PT, T);
	and(P[31], X1[31], X2[9]);
	and(P[30], X1[30], X2[9]);
	and(P[29], X1[29], X2[9]);
	and(P[28], X1[28], X2[9]);
	and(P[27], X1[27], X2[9]);
	and(P[26], X1[26], X2[9]);
	and(P[25], X1[25], X2[9]);
	and(P[24], X1[24], X2[9]);
	and(P[23], X1[23], X2[9]);
	and(P[22], X1[22], X2[9]);
	and(P[21], X1[21], X2[9]);
	and(P[20], X1[20], X2[9]);
	and(P[19], X1[19], X2[9]);
	and(P[18], X1[18], X2[9]);
	and(P[17], X1[17], X2[9]);
	and(P[16], X1[16], X2[9]);
	and(P[15], X1[15], X2[9]);
	and(P[14], X1[14], X2[9]);
	and(P[13], X1[13], X2[9]);
	and(P[12], X1[12], X2[9]);
	and(P[11], X1[11], X2[9]);
	and(P[10], X1[10], X2[9]);
	and(P[9], X1[9], X2[9]);
	and(P[8], X1[8], X2[9]);
	and(P[7], X1[7], X2[9]);
	and(P[6], X1[6], X2[9]);
	and(P[5], X1[5], X2[9]);
	and(P[4], X1[4], X2[9]);
	and(P[3], X1[3], X2[9]);
	and(P[2], X1[2], X2[9]);
	and(P[1], X1[1], X2[9]);
	and(P[0], X1[0], X2[9]);
	fulladd fadd9 (T, PT, P);
	leftmove lm9 (PT, T);
	and(P[31], X1[31], X2[8]);
	and(P[30], X1[30], X2[8]);
	and(P[29], X1[29], X2[8]);
	and(P[28], X1[28], X2[8]);
	and(P[27], X1[27], X2[8]);
	and(P[26], X1[26], X2[8]);
	and(P[25], X1[25], X2[8]);
	and(P[24], X1[24], X2[8]);
	and(P[23], X1[23], X2[8]);
	and(P[22], X1[22], X2[8]);
	and(P[21], X1[21], X2[8]);
	and(P[20], X1[20], X2[8]);
	and(P[19], X1[19], X2[8]);
	and(P[18], X1[18], X2[8]);
	and(P[17], X1[17], X2[8]);
	and(P[16], X1[16], X2[8]);
	and(P[15], X1[15], X2[8]);
	and(P[14], X1[14], X2[8]);
	and(P[13], X1[13], X2[8]);
	and(P[12], X1[12], X2[8]);
	and(P[11], X1[11], X2[8]);
	and(P[10], X1[10], X2[8]);
	and(P[9], X1[9], X2[8]);
	and(P[8], X1[8], X2[8]);
	and(P[7], X1[7], X2[8]);
	and(P[6], X1[6], X2[8]);
	and(P[5], X1[5], X2[8]);
	and(P[4], X1[4], X2[8]);
	and(P[3], X1[3], X2[8]);
	and(P[2], X1[2], X2[8]);
	and(P[1], X1[1], X2[8]);
	and(P[0], X1[0], X2[8]);
	fulladd fadd8 (T, PT, P);
	leftmove lm8 (PT, T);
	and(P[31], X1[31], X2[7]);
	and(P[30], X1[30], X2[7]);
	and(P[29], X1[29], X2[7]);
	and(P[28], X1[28], X2[7]);
	and(P[27], X1[27], X2[7]);
	and(P[26], X1[26], X2[7]);
	and(P[25], X1[25], X2[7]);
	and(P[24], X1[24], X2[7]);
	and(P[23], X1[23], X2[7]);
	and(P[22], X1[22], X2[7]);
	and(P[21], X1[21], X2[7]);
	and(P[20], X1[20], X2[7]);
	and(P[19], X1[19], X2[7]);
	and(P[18], X1[18], X2[7]);
	and(P[17], X1[17], X2[7]);
	and(P[16], X1[16], X2[7]);
	and(P[15], X1[15], X2[7]);
	and(P[14], X1[14], X2[7]);
	and(P[13], X1[13], X2[7]);
	and(P[12], X1[12], X2[7]);
	and(P[11], X1[11], X2[7]);
	and(P[10], X1[10], X2[7]);
	and(P[9], X1[9], X2[7]);
	and(P[8], X1[8], X2[7]);
	and(P[7], X1[7], X2[7]);
	and(P[6], X1[6], X2[7]);
	and(P[5], X1[5], X2[7]);
	and(P[4], X1[4], X2[7]);
	and(P[3], X1[3], X2[7]);
	and(P[2], X1[2], X2[7]);
	and(P[1], X1[1], X2[7]);
	and(P[0], X1[0], X2[7]);
	fulladd fadd7 (T, PT, P);
	leftmove lm7 (PT, T);
	and(P[31], X1[31], X2[6]);
	and(P[30], X1[30], X2[6]);
	and(P[29], X1[29], X2[6]);
	and(P[28], X1[28], X2[6]);
	and(P[27], X1[27], X2[6]);
	and(P[26], X1[26], X2[6]);
	and(P[25], X1[25], X2[6]);
	and(P[24], X1[24], X2[6]);
	and(P[23], X1[23], X2[6]);
	and(P[22], X1[22], X2[6]);
	and(P[21], X1[21], X2[6]);
	and(P[20], X1[20], X2[6]);
	and(P[19], X1[19], X2[6]);
	and(P[18], X1[18], X2[6]);
	and(P[17], X1[17], X2[6]);
	and(P[16], X1[16], X2[6]);
	and(P[15], X1[15], X2[6]);
	and(P[14], X1[14], X2[6]);
	and(P[13], X1[13], X2[6]);
	and(P[12], X1[12], X2[6]);
	and(P[11], X1[11], X2[6]);
	and(P[10], X1[10], X2[6]);
	and(P[9], X1[9], X2[6]);
	and(P[8], X1[8], X2[6]);
	and(P[7], X1[7], X2[6]);
	and(P[6], X1[6], X2[6]);
	and(P[5], X1[5], X2[6]);
	and(P[4], X1[4], X2[6]);
	and(P[3], X1[3], X2[6]);
	and(P[2], X1[2], X2[6]);
	and(P[1], X1[1], X2[6]);
	and(P[0], X1[0], X2[6]);
	fulladd fadd6 (T, PT, P);
	leftmove lm6 (PT, T);
	and(P[31], X1[31], X2[5]);
	and(P[30], X1[30], X2[5]);
	and(P[29], X1[29], X2[5]);
	and(P[28], X1[28], X2[5]);
	and(P[27], X1[27], X2[5]);
	and(P[26], X1[26], X2[5]);
	and(P[25], X1[25], X2[5]);
	and(P[24], X1[24], X2[5]);
	and(P[23], X1[23], X2[5]);
	and(P[22], X1[22], X2[5]);
	and(P[21], X1[21], X2[5]);
	and(P[20], X1[20], X2[5]);
	and(P[19], X1[19], X2[5]);
	and(P[18], X1[18], X2[5]);
	and(P[17], X1[17], X2[5]);
	and(P[16], X1[16], X2[5]);
	and(P[15], X1[15], X2[5]);
	and(P[14], X1[14], X2[5]);
	and(P[13], X1[13], X2[5]);
	and(P[12], X1[12], X2[5]);
	and(P[11], X1[11], X2[5]);
	and(P[10], X1[10], X2[5]);
	and(P[9], X1[9], X2[5]);
	and(P[8], X1[8], X2[5]);
	and(P[7], X1[7], X2[5]);
	and(P[6], X1[6], X2[5]);
	and(P[5], X1[5], X2[5]);
	and(P[4], X1[4], X2[5]);
	and(P[3], X1[3], X2[5]);
	and(P[2], X1[2], X2[5]);
	and(P[1], X1[1], X2[5]);
	and(P[0], X1[0], X2[5]);
	fulladd fadd5 (T, PT, P);
	leftmove lm5 (PT, T);
	and(P[31], X1[31], X2[4]);
	and(P[30], X1[30], X2[4]);
	and(P[29], X1[29], X2[4]);
	and(P[28], X1[28], X2[4]);
	and(P[27], X1[27], X2[4]);
	and(P[26], X1[26], X2[4]);
	and(P[25], X1[25], X2[4]);
	and(P[24], X1[24], X2[4]);
	and(P[23], X1[23], X2[4]);
	and(P[22], X1[22], X2[4]);
	and(P[21], X1[21], X2[4]);
	and(P[20], X1[20], X2[4]);
	and(P[19], X1[19], X2[4]);
	and(P[18], X1[18], X2[4]);
	and(P[17], X1[17], X2[4]);
	and(P[16], X1[16], X2[4]);
	and(P[15], X1[15], X2[4]);
	and(P[14], X1[14], X2[4]);
	and(P[13], X1[13], X2[4]);
	and(P[12], X1[12], X2[4]);
	and(P[11], X1[11], X2[4]);
	and(P[10], X1[10], X2[4]);
	and(P[9], X1[9], X2[4]);
	and(P[8], X1[8], X2[4]);
	and(P[7], X1[7], X2[4]);
	and(P[6], X1[6], X2[4]);
	and(P[5], X1[5], X2[4]);
	and(P[4], X1[4], X2[4]);
	and(P[3], X1[3], X2[4]);
	and(P[2], X1[2], X2[4]);
	and(P[1], X1[1], X2[4]);
	and(P[0], X1[0], X2[4]);
	fulladd fadd4 (T, PT, P);
	leftmove lm4 (PT, T);
	and(P[31], X1[31], X2[3]);
	and(P[30], X1[30], X2[3]);
	and(P[29], X1[29], X2[3]);
	and(P[28], X1[28], X2[3]);
	and(P[27], X1[27], X2[3]);
	and(P[26], X1[26], X2[3]);
	and(P[25], X1[25], X2[3]);
	and(P[24], X1[24], X2[3]);
	and(P[23], X1[23], X2[3]);
	and(P[22], X1[22], X2[3]);
	and(P[21], X1[21], X2[3]);
	and(P[20], X1[20], X2[3]);
	and(P[19], X1[19], X2[3]);
	and(P[18], X1[18], X2[3]);
	and(P[17], X1[17], X2[3]);
	and(P[16], X1[16], X2[3]);
	and(P[15], X1[15], X2[3]);
	and(P[14], X1[14], X2[3]);
	and(P[13], X1[13], X2[3]);
	and(P[12], X1[12], X2[3]);
	and(P[11], X1[11], X2[3]);
	and(P[10], X1[10], X2[3]);
	and(P[9], X1[9], X2[3]);
	and(P[8], X1[8], X2[3]);
	and(P[7], X1[7], X2[3]);
	and(P[6], X1[6], X2[3]);
	and(P[5], X1[5], X2[3]);
	and(P[4], X1[4], X2[3]);
	and(P[3], X1[3], X2[3]);
	and(P[2], X1[2], X2[3]);
	and(P[1], X1[1], X2[3]);
	and(P[0], X1[0], X2[3]);
	fulladd fadd3 (T, PT, P);
	leftmove lm3 (PT, T);
	and(P[31], X1[31], X2[2]);
	and(P[30], X1[30], X2[2]);
	and(P[29], X1[29], X2[2]);
	and(P[28], X1[28], X2[2]);
	and(P[27], X1[27], X2[2]);
	and(P[26], X1[26], X2[2]);
	and(P[25], X1[25], X2[2]);
	and(P[24], X1[24], X2[2]);
	and(P[23], X1[23], X2[2]);
	and(P[22], X1[22], X2[2]);
	and(P[21], X1[21], X2[2]);
	and(P[20], X1[20], X2[2]);
	and(P[19], X1[19], X2[2]);
	and(P[18], X1[18], X2[2]);
	and(P[17], X1[17], X2[2]);
	and(P[16], X1[16], X2[2]);
	and(P[15], X1[15], X2[2]);
	and(P[14], X1[14], X2[2]);
	and(P[13], X1[13], X2[2]);
	and(P[12], X1[12], X2[2]);
	and(P[11], X1[11], X2[2]);
	and(P[10], X1[10], X2[2]);
	and(P[9], X1[9], X2[2]);
	and(P[8], X1[8], X2[2]);
	and(P[7], X1[7], X2[2]);
	and(P[6], X1[6], X2[2]);
	and(P[5], X1[5], X2[2]);
	and(P[4], X1[4], X2[2]);
	and(P[3], X1[3], X2[2]);
	and(P[2], X1[2], X2[2]);
	and(P[1], X1[1], X2[2]);
	and(P[0], X1[0], X2[2]);
	fulladd fadd2 (T, PT, P);
	leftmove lm2 (PT, T);
	and(P[31], X1[31], X2[1]);
	and(P[30], X1[30], X2[1]);
	and(P[29], X1[29], X2[1]);
	and(P[28], X1[28], X2[1]);
	and(P[27], X1[27], X2[1]);
	and(P[26], X1[26], X2[1]);
	and(P[25], X1[25], X2[1]);
	and(P[24], X1[24], X2[1]);
	and(P[23], X1[23], X2[1]);
	and(P[22], X1[22], X2[1]);
	and(P[21], X1[21], X2[1]);
	and(P[20], X1[20], X2[1]);
	and(P[19], X1[19], X2[1]);
	and(P[18], X1[18], X2[1]);
	and(P[17], X1[17], X2[1]);
	and(P[16], X1[16], X2[1]);
	and(P[15], X1[15], X2[1]);
	and(P[14], X1[14], X2[1]);
	and(P[13], X1[13], X2[1]);
	and(P[12], X1[12], X2[1]);
	and(P[11], X1[11], X2[1]);
	and(P[10], X1[10], X2[1]);
	and(P[9], X1[9], X2[1]);
	and(P[8], X1[8], X2[1]);
	and(P[7], X1[7], X2[1]);
	and(P[6], X1[6], X2[1]);
	and(P[5], X1[5], X2[1]);
	and(P[4], X1[4], X2[1]);
	and(P[3], X1[3], X2[1]);
	and(P[2], X1[2], X2[1]);
	and(P[1], X1[1], X2[1]);
	and(P[0], X1[0], X2[1]);
	fulladd fadd1 (T, PT, P);
	leftmove lm1 (PT, T);
	and(P[31], X1[31], X2[0]);
	and(P[30], X1[30], X2[0]);
	and(P[29], X1[29], X2[0]);
	and(P[28], X1[28], X2[0]);
	and(P[27], X1[27], X2[0]);
	and(P[26], X1[26], X2[0]);
	and(P[25], X1[25], X2[0]);
	and(P[24], X1[24], X2[0]);
	and(P[23], X1[23], X2[0]);
	and(P[22], X1[22], X2[0]);
	and(P[21], X1[21], X2[0]);
	and(P[20], X1[20], X2[0]);
	and(P[19], X1[19], X2[0]);
	and(P[18], X1[18], X2[0]);
	and(P[17], X1[17], X2[0]);
	and(P[16], X1[16], X2[0]);
	and(P[15], X1[15], X2[0]);
	and(P[14], X1[14], X2[0]);
	and(P[13], X1[13], X2[0]);
	and(P[12], X1[12], X2[0]);
	and(P[11], X1[11], X2[0]);
	and(P[10], X1[10], X2[0]);
	and(P[9], X1[9], X2[0]);
	and(P[8], X1[8], X2[0]);
	and(P[7], X1[7], X2[0]);
	and(P[6], X1[6], X2[0]);
	and(P[5], X1[5], X2[0]);
	and(P[4], X1[4], X2[0]);
	and(P[3], X1[3], X2[0]);
	and(P[2], X1[2], X2[0]);
	and(P[1], X1[1], X2[0]);
	and(P[0], X1[0], X2[0]);
	fulladd fadd0 (T, PT, P);
	leftmove lm0 (PT, T);
	buf(F[31], T[31]);
	buf(F[30], T[30]);
	buf(F[29], T[29]);
	buf(F[28], T[28]);
	buf(F[27], T[27]);
	buf(F[26], T[26]);
	buf(F[25], T[25]);
	buf(F[24], T[24]);
	buf(F[23], T[23]);
	buf(F[22], T[22]);
	buf(F[21], T[21]);
	buf(F[20], T[20]);
	buf(F[19], T[19]);
	buf(F[18], T[18]);
	buf(F[17], T[17]);
	buf(F[16], T[16]);
	buf(F[15], T[15]);
	buf(F[14], T[14]);
	buf(F[13], T[13]);
	buf(F[12], T[12]);
	buf(F[11], T[11]);
	buf(F[10], T[10]);
	buf(F[9], T[9]);
	buf(F[8], T[8]);
	buf(F[7], T[7]);
	buf(F[6], T[6]);
	buf(F[5], T[5]);
	buf(F[4], T[4]);
	buf(F[3], T[3]);
	buf(F[2], T[2]);
	buf(F[1], T[1]);
	buf(F[0], T[0]);
	
endmodule
